module module7SEG(
    input logic [3:0] cod_bin;
    output logic [1:0] anodo_po;
    output logic [6:0] catodo_po;
)

    assign A = cod_bin[3];
    assign B = cod_bin[2];
    assign C = cod_bin[1];
    assign D = cod_bin[0];

    //seg a
    assign seg_a = ;
    
    //seg b
    //seg c
    //seg d
    //seg e
    //seg f
    //seg g

endmodule